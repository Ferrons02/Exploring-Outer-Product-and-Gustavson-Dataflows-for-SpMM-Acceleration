/usr/pack/gf-22-kgf/dz/openroad/10M_2Mx_6Cx_2Ix_LB__PLUS-V1.0_3.0a/22FDSOI_10M_2Mx_6Cx_2Ix_LB_104cpp_6p75t_openaroad_tech.lef