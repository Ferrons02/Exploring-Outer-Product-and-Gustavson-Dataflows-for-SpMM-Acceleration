/usr/pack/gf-22-kgf/dz/innovus/10M_2Mx_6Cx_2Ix_LB__PLUS-V1.0_3.0a/22FDSOI_10M_2Mx_6Cx_2Ix_LB_104cpp_tech.lef