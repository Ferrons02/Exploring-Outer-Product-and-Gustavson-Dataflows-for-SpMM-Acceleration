/usr/pack/gf-22-kgf/invecas/io/2020.01/IN22FDX_GPIO18_10M3S40PI_FE_RELV02R02SZ/lef.dz/IN22FDX_GPIO18_10M3S40PI.lef