/usr/pack/gf-22-kgf/invecas/std8t/2020.01/GF22FDX_SC8T_104CPP_BASE_CSC28SL_FDK_RELV06R40/lef/GF22FDX_SC8T_104CPP_BASE_CSC28SL.lef